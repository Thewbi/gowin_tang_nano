// the state machine that runs the demo application has three states: IDLE, SEND and WAIT
//
// IDLE is entered on reset. IDLE immediately transitions to SEND.
// IDLE does not perform any action.
//
// SEND is entered after IDLE and when the wait period is over.
// During SEND a string of DATA_NUM characters is transmitted, one
// character per clock tick. Once all characters are transmitted,
// the transition to WAIT takes place because the demo wants to 
// wait around for some time before sending DATA_NUM characters again.
//
// In WAIT, the system remains still whithout sending data for one
// second. WAIT is the only state, where the system checks for incoming data.
// If a byte is received, that exact byte is immediately sent out over the tx line.
// 

module top(

    // input
    input wire sys_clk,         // clk input
    input wire sys_rst_n,       // reset input button  (active low)
	input wire uart_rx,         // UART RX
    input wire btn1_n,          // push button 1 (active low)
    input wire jtag_clk,
    input wire jtag_tdi,
    input wire jtag_tms,

    // output
    output wire [5:0] led,      // 6 LEDS pin
	output wire uart_tx,        // UART TX
    output wire jtag_tdo

);


/**/
//
// wishbone
//

wire [31:0] read_data;
wire [31:0] write_data;
wire ack;
wire cyc;
wire stb;
wire [31:0] addr;
wire we;

wire start_read_transaction; // output by the JTAG tap to cause the withbone master to read the slave
wire start_write_transaction; // output by the JTAG tap to cause the withbone master to write the slave
wire[7:0] wishbone_tx_data;

wishbone_master wb_master (

    // input
    .clk_i(sys_clk),
    .rst_i(~sys_rst_n),

    // input master
    .data_i(read_data),
    .ack_i(ack),

    // input wbi custom 
    .start_read_transaction_i(start_read_transaction),
    .start_write_transaction_i(start_write_transaction),
    .write_transaction_data_i(wishbone_tx_data),
    
    // output master
    .addr_o(addr),
    .we_o(we),
    .data_o(write_data), // output to the slave on write transactions
    .cyc_o(cyc),
    .stb_o(stb),

    // output wbi custom
    .read_transaction_data_o()

);



//
// Timer - perform action every second
//

parameter BAUD_RATE = 115200; // serial baud rate, 115200 bits per second
parameter CLK_FRE_MHZ = CLK_FRE * 1000000;
parameter CYCLES_PER_BIT = CLK_FRE_MHZ / BAUD_RATE; // CLOCK TICKS per bit

/*
reg [31:0] counter;
reg [7:0] tx_counter;

always @(posedge sys_clk)
begin
    counter = counter + 1;

    if (counter == CLK_FRE_MHZ)
    begin

        counter = 32'd0;

        // perform action every second

// Enable this snippet for the wishbone RX slave
//        // start/stop a wishbone read transaction
//        start_read_transaction <= ~start_read_transaction;
//

//        // start the wishbone write transaction
//        start_write_transaction = 1;
//        tx_data = tx_data + 1;

//        // transmit data over the raw UART TX (without wishbone)
//        tx_data_valid = ~tx_data_valid;
//        tx_data = 8'h01;

    end

//    // ENABLE this for UART TX write
//    if (counter >= (CYCLES_PER_BIT * 8))
//    begin
//        // stop the wishbone write transaction
//        start_write_transaction = 0;
//    end

end
*/




//
// UART demo application
//

//
// combinational logic for UART
//

parameter DATA_NUM = 22;
wire [DATA_NUM * 8 - 1:0] send_data;
// DEBUG control the uart tx
//reg printf = 1'b0;
wire printf;

reg[7:0]                        tx_str;

wire[7:0]                       tx_data;
wire[7:0]                       tx_cnt;

wire                            tx_data_ready; // output of the tx module. Asserted when transmission has been performed
wire[7:0]                       rx_data;
reg                             rx_data_ready = 1'b1; // receiving data is always enabled
wire                            tx_data_valid;

uart_controller 
#(
    .DATA_NUM(DATA_NUM)
) uart_controller_inst (

    // input
	.clk                        (sys_clk),
	.rst_n                      (sys_rst_n),
    .tx_str                     (tx_str),
    .printf                     (printf),
    .tx_data_ready              (tx_data_ready),
    .o_tx_data_valid            (tx_data_valid),
    .rx_data                    (rx_data),
    .rx_data_valid              (rx_data_valid),

    // output
    .o_tx_cnt                   (tx_cnt),
	.o_tx_data                  (tx_data)
    
);

parameter                        CLK_FRE  = 27; // Mhz. The Tang Nano 9K has a 27 Mhz clock source on board
parameter                        UART_FRE = 115200; // baudrate

always @(*)
begin
	tx_str <= send_data[(DATA_NUM - 1 - tx_cnt) * 8 +: 8];
end

uart_rx
#(
	.CLK_FRE(CLK_FRE),
	.BAUD_RATE(UART_FRE)
) uart_rx_inst (
    // input
	.clk                        (sys_clk),
	.rst_n                      (sys_rst_n),	
	.rx_data_ready              (rx_data_ready),
	.rx_pin                     (uart_rx),

    // output
    .rx_data                    (rx_data),
	.rx_data_valid              (rx_data_valid)
);

uart_tx
#(
	.CLK_FRE(CLK_FRE),
	.BAUD_RATE(UART_FRE)
) uart_tx_inst (
    // input
	.clk                        (sys_clk),
	.rst_n                      (sys_rst_n),
	.tx_data                    (tx_data),
	.tx_data_valid              (tx_data_valid),

    // output
	.tx_data_ready              (tx_data_ready),
	.tx_pin                     (uart_tx)
);

//
// user button demo application
//

// http://nandland.com/project-4-debounce-a-switch/

reg  r_Switch_1 = 1'b0;
wire w_Switch_1;

// Instantiate Debounce Module
Debounce_Switch debounce_Inst
(
    .i_Clk(sys_clk), 
    .i_Switch(btn1_n),
    .o_Switch(w_Switch_1)
);


//
// JTAG example
//

reg r_LED_1 = 1'b0;
wire [5:0] leds;
reg [5:0] r_led_reg = 6'b111111;

always @(leds)
begin
    r_led_reg <= leds;
end

jtag_tap #(
    .DATA_NUM(DATA_NUM)
) jtag_tap_inst (

    //
    // JTAG
    //

    // input
    .clk(sys_clk),
    .rst_n(sys_rst_n),
    .jtag_clk(jtag_clk),
    .jtag_tdi(jtag_tdi),
    .jtag_tms(jtag_tms),
    
    // output    
    .jtag_tdo(jtag_tdo),

    // debug output
    .r_led_reg(leds),

    // printf output enabled
    .send_data(send_data),
    .printf(printf),

    // printf output disabled
    //.send_data(),
    //.printf(),

    // when a JTAG command for dmi (0x11) arrives, the JTAG_TAP will
    // output commands to the wishbone master here. The wishbone master
    // talks to the RISCV DM which is a wishbone slave.
    .start_read_transaction_o(start_read_transaction),
    .start_write_transaction_o(start_write_transaction),
    .write_transaction_data_o(wishbone_tx_data)

);

//
// wishbone
//

wishbone_led_slave #(
    .DATA_NUM(DATA_NUM)
) wb_led_slave (

    // input
    .clk_i(sys_clk),
    .rst_i(~sys_rst_n),

    // input slave
    .addr_i(addr), // address within a wishbone slave
    .we_i(we),
    .data_i(write_data), // the master places the data to write into write_data
    .cyc_i(cyc),
    .stb_i(stb),

    // input custom

    // output slave
    .data_o(read_data), // the TX slave does not use data_o. It does not return any usefull data.
    .ack_o(ack),

    // output wbi
    .led_port_o(led) // output to the LEDs port

    // printf - does not work because it causes a logical cycle, the state machine is not clocked
    //.send_data(send_data),
    //.printf(printf)

);

endmodule