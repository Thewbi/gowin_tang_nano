//module top (
//    input sys_clk,          // clk input
//    input sys_rst_n,        // reset input
//    output reg [5:0] led    // 6 LEDS pin
//);

//reg [23:0] counter;

// // update the counter variable
//always @(posedge sys_clk or negedge sys_rst_n) begin
//    if (!sys_rst_n)
//        counter <= 24'd0;
//    else if (counter < 24'd1349_9999)       // 0.5s delay
//        counter <= counter + 1'b1;
//    else
//        counter <= 24'd0;
//end


// // update the LEDs
//always @(posedge sys_clk or negedge sys_rst_n) begin
//    if (!sys_rst_n)
//        led <= 6'b111110;
//    else if (counter == 24'd1349_9999)       // 0.5s delay
//        led[5:0] <= {led[4:0],led[5]};    // left to right
//        led[5:0] <= {led[0], led[5:1]};     // right to left
//    else
//        led <= led;
//end

//endmodule